
module system (
	clk_clk,
	sw_wire_export,
	led_wire_leds);	

	input		clk_clk;
	input	[9:0]	sw_wire_export;
	output	[9:0]	led_wire_leds;
endmodule
